`timescale 1 ns / 1 ps

module axi_cfg_register #
(
